** Profile: "SCHEMATIC1-OpAmpSim"  [ Z:\Tim File Sync\work\HandTie\HandTieCode\OrCAD\HandTieHardwareSim\handtiesimulation2-pspicefiles\schematic1\opampsim.sim ] 

** Creating circuit file "OpAmpSim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/OrCAD/OrCAD_16.5_Lite/tools/capture/library/CustomLibrary/LM6132B.lib" 
.LIB "C:/OrCAD/OrCAD_16.5_Lite/tools/capture/library/CustomLibrary/LM6132A.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
